CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
120 130 30 80 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
56
13 Logic Switch~
5 234 336 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 29424 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9840 0 0
2
43087.6 7
0
13 Logic Switch~
5 233 414 0 1 11
0 11
0
0 0 29424 0
2 0V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6910 0 0
2
43087.6 6
0
13 Logic Switch~
5 217 560 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 29424 0
2 5V
-6 -16 8 -8
2 RD
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
449 0 0
2
43087.6 5
0
13 Logic Switch~
5 215 606 0 10 11
0 41 0 0 0 0 0 0 0 0
1
0
0 0 29424 0
2 5V
-6 -16 8 -8
2 CS
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8761 0 0
2
43087.6 4
0
13 Logic Switch~
5 214 648 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 29424 0
2 5V
-6 -16 8 -8
2 OE
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6748 0 0
2
43087.6 3
0
13 Logic Switch~
5 593 203 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 I0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7393 0 0
2
43087.6 2
0
13 Logic Switch~
5 720 195 0 10 11
0 30 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 I1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7699 0 0
2
43087.6 1
0
13 Logic Switch~
5 830 191 0 1 11
0 29
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 I2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6638 0 0
2
43087.6 0
0
9 2-In AND~
219 358 427 0 3 22
0 10 2 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
4595 0 0
2
43087.6 0
0
9 2-In AND~
219 358 376 0 3 22
0 12 11 5
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U37D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
9395 0 0
2
43087.6 0
0
9 Inverter~
13 280 316 0 2 22
0 10 12
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U24C
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 24 0
1 U
3303 0 0
2
43087.6 53
0
9 Inverter~
13 280 383 0 2 22
0 11 2
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U24D
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 24 0
1 U
4498 0 0
2
43087.6 52
0
9 2-In AND~
219 359 324 0 3 22
0 12 2 7
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U22C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 22 0
1 U
9728 0 0
2
43087.6 51
0
7 Pulser~
4 202 499 0 10 12
0 46 47 48 45 0 0 5 5 1
8
0
0 0 4144 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3789 0 0
2
43087.6 50
0
5 7415~
219 324 525 0 4 22
0 45 44 41 9
0
0 0 112 0
6 74LS15
-21 -28 21 -20
4 U15C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 20 0
1 U
3978 0 0
2
43087.6 49
0
5 7415~
219 371 639 0 4 22
0 42 41 43 16
0
0 0 112 0
6 74LS15
-21 -28 21 -20
4 U25A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 25 0
1 U
3494 0 0
2
43087.6 48
0
9 Inverter~
13 270 525 0 2 22
0 42 44
0
0 0 112 0
6 74LS04
-21 -19 21 -11
4 U24E
-14 -20 14 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 24 0
1 U
3507 0 0
2
43087.6 47
0
9 2-In AND~
219 475 333 0 3 22
0 7 9 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U22D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 22 0
1 U
5151 0 0
2
43087.6 46
0
9 2-In AND~
219 474 385 0 3 22
0 5 9 6
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U26A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 26 0
1 U
3701 0 0
2
43087.6 45
0
9 2-In AND~
219 474 436 0 3 22
0 3 9 4
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U26B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 26 0
1 U
8585 0 0
2
43087.6 44
0
12 D Flip-Flop~
219 655 328 0 4 9
0 31 8 49 40
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U27
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8809 0 0
2
43087.6 43
0
12 D Flip-Flop~
219 767 328 0 4 9
0 30 8 50 39
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U28
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5993 0 0
2
43087.6 42
0
12 D Flip-Flop~
219 869 328 0 4 9
0 29 8 51 38
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U29
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8654 0 0
2
43087.6 41
0
9 2-In AND~
219 705 371 0 3 22
0 40 7 32
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U26C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 26 0
1 U
7223 0 0
2
43087.6 40
0
9 2-In AND~
219 811 370 0 3 22
0 39 7 23
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U26D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 26 0
1 U
3641 0 0
2
43087.6 39
0
9 2-In AND~
219 934 369 0 3 22
0 38 7 20
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U30A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 27 0
1 U
3104 0 0
2
43087.6 38
0
14 Logic Display~
6 698 274 0 1 2
10 40
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 I8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3296 0 0
2
43087.6 37
0
14 Logic Display~
6 809 274 0 1 2
10 39
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 I9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8534 0 0
2
43087.6 36
0
14 Logic Display~
6 931 274 0 1 2
10 38
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
949 0 0
2
43087.6 35
0
12 D Flip-Flop~
219 655 466 0 4 9
0 31 6 52 37
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U31
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3371 0 0
2
43087.6 34
0
12 D Flip-Flop~
219 766 464 0 4 9
0 30 6 53 36
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U32
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7311 0 0
2
43087.6 33
0
12 D Flip-Flop~
219 871 462 0 4 9
0 29 6 54 35
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U33
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
43087.6 32
0
9 2-In AND~
219 681 516 0 3 22
0 37 5 33
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U30B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 27 0
1 U
3526 0 0
2
43087.6 31
0
9 2-In AND~
219 794 515 0 3 22
0 36 5 24
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U30C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 27 0
1 U
4129 0 0
2
43087.6 30
0
9 2-In AND~
219 905 514 0 3 22
0 35 5 21
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U30D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 27 0
1 U
6278 0 0
2
43087.6 29
0
14 Logic Display~
6 681 412 0 1 2
10 37
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
43087.6 28
0
14 Logic Display~
6 793 411 0 1 2
10 36
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8323 0 0
2
43087.6 27
0
14 Logic Display~
6 902 409 0 1 2
10 35
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3984 0 0
2
43087.6 26
0
12 D Flip-Flop~
219 636 615 0 4 9
0 31 4 55 28
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U34
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7622 0 0
2
43087.6 25
0
12 D Flip-Flop~
219 751 619 0 4 9
0 30 4 56 27
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U35
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
816 0 0
2
43087.6 24
0
12 D Flip-Flop~
219 856 614 0 4 9
0 29 4 57 26
0
0 0 4208 0
3 DFF
-10 -53 11 -45
3 U36
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4656 0 0
2
43087.6 23
0
9 2-In AND~
219 663 666 0 3 22
0 28 3 34
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U37A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 28 0
1 U
6356 0 0
2
43087.6 22
0
9 2-In AND~
219 776 665 0 3 22
0 27 3 25
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U37B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 28 0
1 U
7479 0 0
2
43087.6 21
0
9 2-In AND~
219 887 663 0 3 22
0 26 3 22
0
0 0 112 270
6 74LS08
-21 -24 21 -16
4 U37C
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 28 0
1 U
5690 0 0
2
43087.6 20
0
8 3-In OR~
219 667 755 0 4 22
0 32 33 34 19
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U11B
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 16 0
1 U
5617 0 0
2
43087.6 19
0
14 Logic Display~
6 666 561 0 1 2
10 28
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3903 0 0
2
43087.6 18
0
14 Logic Display~
6 778 565 0 1 2
10 27
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4452 0 0
2
43087.6 17
0
14 Logic Display~
6 888 560 0 1 2
10 26
0
0 0 53344 0
6 100MEG
3 -16 45 -8
3 I16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6282 0 0
2
43087.6 16
0
8 3-In OR~
219 780 752 0 4 22
0 23 24 25 18
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U11C
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 16 0
1 U
7187 0 0
2
43087.6 15
0
8 3-In OR~
219 891 753 0 4 22
0 20 21 22 17
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U38A
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 29 0
1 U
6866 0 0
2
43087.6 14
0
10 Buffer 3S~
219 895 823 0 3 22
0 17 16 13
0
0 0 624 270
8 BUFFER3S
-27 -51 29 -43
2 D2
21 -5 35 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 12 13 11 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 23 0
1 U
7670 0 0
2
43087.6 13
0
10 Buffer 3S~
219 784 823 0 3 22
0 18 16 14
0
0 0 624 270
8 BUFFER3S
-27 -51 29 -43
2 D1
21 -5 35 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 2 1 3 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
951 0 0
2
43087.6 12
0
10 Buffer 3S~
219 671 822 0 3 22
0 19 16 15
0
0 0 624 270
8 BUFFER3S
-27 -51 29 -43
2 D0
21 -5 35 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
0
22

0 5 4 6 2 1 3 5 4 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
9536 0 0
2
43087.6 11
0
14 Logic Display~
6 670 850 0 1 2
10 15
0
0 0 53344 180
6 100MEG
3 -16 45 -8
3 I17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5495 0 0
2
43087.6 10
0
14 Logic Display~
6 783 852 0 1 2
10 14
0
0 0 53344 180
6 100MEG
3 -16 45 -8
3 I18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8152 0 0
2
43087.6 9
0
14 Logic Display~
6 894 852 0 1 2
10 13
0
0 0 53344 180
6 100MEG
3 -16 45 -8
3 I19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6223 0 0
2
43087.6 8
0
84
2 2 2 0 0 4224 0 12 9 0 0 3
301 383
301 436
334 436
2 0 3 0 0 4096 0 42 0 0 4 2
652 644
652 625
2 0 3 0 0 0 0 43 0 0 4 2
765 643
765 625
0 2 3 0 0 8320 0 0 44 23 0 4
426 427
426 625
876 625
876 641
0 2 4 0 0 4096 0 0 39 7 0 3
601 613
601 597
612 597
0 2 4 0 0 0 0 0 40 7 0 3
718 613
718 601
727 601
3 2 4 0 0 8320 0 20 41 0 0 5
495 436
495 613
825 613
825 596
832 596
2 0 5 0 0 4096 0 33 0 0 10 2
670 494
670 484
2 0 5 0 0 0 0 34 0 0 10 2
783 493
783 484
0 2 5 0 0 8320 0 0 35 24 0 4
409 376
409 484
894 484
894 492
0 2 6 0 0 4096 0 0 30 13 0 3
623 465
623 448
631 448
0 2 6 0 0 4096 0 0 31 13 0 3
736 465
736 446
742 446
3 2 6 0 0 12416 0 19 32 0 0 6
495 385
570 385
570 465
842 465
842 444
847 444
2 0 7 0 0 4096 0 24 0 0 16 2
694 349
694 340
2 0 7 0 0 0 0 25 0 0 16 2
800 348
800 340
0 2 7 0 0 16512 0 0 26 25 0 6
408 324
408 361
653 361
653 340
923 340
923 347
0 2 8 0 0 4096 0 0 21 19 0 3
621 333
621 310
631 310
0 2 8 0 0 0 0 0 22 19 0 3
738 333
738 310
743 310
3 2 8 0 0 4224 0 18 23 0 0 4
496 333
841 333
841 310
845 310
2 0 9 0 0 4096 0 20 0 0 22 2
450 445
433 445
2 0 9 0 0 0 0 19 0 0 22 2
450 394
433 394
4 2 9 0 0 8320 0 15 18 0 0 4
345 525
433 525
433 342
451 342
3 1 3 0 0 0 0 9 20 0 0 2
379 427
450 427
3 1 5 0 0 0 0 10 19 0 0 2
379 376
450 376
3 1 7 0 0 0 0 13 18 0 0 2
380 324
451 324
0 1 10 0 0 4224 0 0 9 84 0 3
257 316
257 418
334 418
1 2 11 0 0 4224 0 2 10 0 0 4
245 414
323 414
323 385
334 385
0 1 12 0 0 4224 0 0 10 30 0 3
323 315
323 367
334 367
2 2 2 0 0 128 0 12 13 0 0 3
301 383
301 333
335 333
2 1 12 0 0 0 0 11 13 0 0 3
301 316
301 315
335 315
1 3 13 0 0 4224 0 56 51 0 0 2
894 838
894 839
1 3 14 0 0 4224 0 55 52 0 0 2
783 838
783 839
1 3 15 0 0 4224 0 54 53 0 0 2
670 836
670 838
0 2 16 0 0 4096 0 0 53 36 0 3
642 797
642 823
659 823
0 2 16 0 0 4096 0 0 52 36 0 3
752 797
752 824
772 824
4 2 16 0 0 8320 0 16 51 0 0 5
392 639
392 797
872 797
872 824
883 824
4 1 17 0 0 4224 0 50 51 0 0 2
894 783
894 809
4 1 18 0 0 4224 0 49 52 0 0 2
783 782
783 809
4 1 19 0 0 4224 0 45 53 0 0 2
670 785
670 808
3 1 20 0 0 4224 0 26 50 0 0 4
932 392
932 723
903 723
903 737
3 2 21 0 0 4224 0 35 50 0 0 4
903 537
903 718
894 718
894 738
3 3 22 0 0 4224 0 50 44 0 0 2
885 737
885 686
3 1 23 0 0 4224 0 25 49 0 0 4
809 393
809 728
792 728
792 736
3 2 24 0 0 4224 0 34 49 0 0 4
792 538
792 722
783 722
783 737
3 3 25 0 0 4224 0 49 43 0 0 2
774 736
774 688
1 0 26 0 0 0 0 48 0 0 61 2
888 578
888 578
1 0 27 0 0 0 0 47 0 0 62 2
778 583
778 583
1 0 28 0 0 0 0 46 0 0 63 2
666 579
666 579
1 0 29 0 0 4096 0 23 0 0 51 2
845 292
832 292
1 0 29 0 0 4096 0 32 0 0 51 2
847 426
832 426
1 1 29 0 0 8320 0 8 41 0 0 3
830 203
832 203
832 578
1 0 30 0 0 4096 0 22 0 0 54 2
743 292
720 292
1 0 30 0 0 0 0 31 0 0 54 2
742 428
720 428
1 1 30 0 0 4224 0 7 40 0 0 3
720 207
720 583
727 583
1 0 31 0 0 4096 0 21 0 0 57 2
631 292
593 292
1 0 31 0 0 0 0 30 0 0 57 2
631 430
593 430
1 1 31 0 0 4224 0 6 39 0 0 3
593 215
593 579
612 579
3 1 32 0 0 4224 0 24 45 0 0 4
703 394
703 718
679 718
679 739
3 2 33 0 0 4224 0 33 45 0 0 4
679 539
679 713
670 713
670 740
3 3 34 0 0 4224 0 42 45 0 0 2
661 689
661 739
4 1 26 0 0 8320 0 41 44 0 0 3
880 578
894 578
894 641
4 1 27 0 0 8320 0 40 43 0 0 3
775 583
783 583
783 643
4 1 28 0 0 8320 0 39 42 0 0 3
660 579
670 579
670 644
1 0 35 0 0 4096 0 38 0 0 67 2
902 427
902 426
1 0 36 0 0 4096 0 37 0 0 68 2
793 429
793 428
1 0 37 0 0 0 0 36 0 0 69 2
681 430
681 430
4 1 35 0 0 8320 0 32 35 0 0 3
895 426
912 426
912 492
4 1 36 0 0 8320 0 31 34 0 0 3
790 428
801 428
801 493
4 1 37 0 0 8320 0 30 33 0 0 3
679 430
688 430
688 494
1 0 38 0 0 0 0 29 0 0 73 2
931 292
931 292
1 0 39 0 0 0 0 28 0 0 74 2
809 292
809 292
1 0 40 0 0 0 0 27 0 0 75 2
698 292
698 292
4 1 38 0 0 8320 0 23 26 0 0 3
893 292
941 292
941 347
4 1 39 0 0 8320 0 22 25 0 0 3
791 292
818 292
818 348
4 1 40 0 0 8320 0 21 24 0 0 3
679 292
712 292
712 349
0 2 41 0 0 8192 0 0 16 77 0 3
292 606
292 639
347 639
1 3 41 0 0 8320 0 4 15 0 0 4
227 606
292 606
292 534
300 534
1 1 42 0 0 8320 0 3 16 0 0 3
229 560
229 630
347 630
1 3 43 0 0 4224 0 5 16 0 0 2
226 648
347 648
1 1 42 0 0 0 0 3 17 0 0 3
229 560
229 525
255 525
2 2 44 0 0 4224 0 17 15 0 0 2
291 525
300 525
4 1 45 0 0 4224 0 14 15 0 0 4
232 499
293 499
293 516
300 516
1 1 11 0 0 0 0 2 12 0 0 3
245 414
245 383
265 383
1 1 10 0 0 0 0 1 11 0 0 3
246 336
246 316
265 316
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
