CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
320 170 30 80 10
176 80 1358 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
16 C:\CM60S\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
0
0
0
0
0
56
13 Logic Switch~
5 853 251 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 Y
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
449 0 0
2
43055.8 15
0
13 Logic Switch~
5 831 251 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 X
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8761 0 0
2
43055.8 14
0
13 Logic Switch~
5 880 252 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 Cin
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6748 0 0
2
43055.8 13
0
13 Logic Switch~
5 654 210 0 1 11
0 50
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 D
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7393 0 0
2
43055.8 3
0
13 Logic Switch~
5 464 211 0 10 11
0 57 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7699 0 0
2
43055.8 4
0
13 Logic Switch~
5 536 212 0 1 11
0 52
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6638 0 0
2
43055.8 5
0
13 Logic Switch~
5 590 212 0 1 11
0 54
0
0 0 21360 270
2 0V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4595 0 0
2
43055.8 6
0
14 Logic Display~
6 1211 414 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 Cout
-15 -21 13 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9395 0 0
2
43055.8 0
0
9 2-In AND~
219 1190 432 0 3 22
0 15 14 3
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U18B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 22 0
1 U
3303 0 0
2
43055.8 0
0
8 2-In OR~
219 1105 401 0 3 22
0 5 7 15
0
0 0 112 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
4498 0 0
2
43055.8 12
0
9 2-In AND~
219 1054 374 0 3 22
0 12 19 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U15A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 19 0
1 U
9728 0 0
2
43055.8 11
0
8 2-In OR~
219 1107 468 0 3 22
0 8 9 14
0
0 0 112 0
6 74LS32
-21 -24 21 -16
4 U12C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3789 0 0
2
43055.8 10
0
9 2-In AND~
219 1040 477 0 3 22
0 6 10 9
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U15B
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 19 0
1 U
3978 0 0
2
43055.8 9
0
8 2-In OR~
219 968 486 0 3 22
0 12 19 10
0
0 0 112 0
6 74LS32
-21 -24 21 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
3494 0 0
2
43055.8 8
0
9 2-In XOR~
219 970 438 0 3 22
0 4 20 6
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 U16A
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
3507 0 0
2
43055.8 7
0
9 2-In AND~
219 914 458 0 3 22
0 7 18 20
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U15C
-17 -24 11 -16
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 19 0
1 U
5151 0 0
2
43055.8 6
0
9 2-In AND~
219 915 413 0 3 22
0 5 11 4
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U15D
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 19 0
1 U
3701 0 0
2
43055.8 5
0
9 Inverter~
13 810 280 0 2 22
0 11 18
0
0 0 112 270
6 74LS04
-21 -19 21 -11
4 U13B
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 17 0
1 U
8585 0 0
2
43055.8 4
0
8 2-In OR~
219 1000 348 0 3 22
0 5 7 21
0
0 0 112 0
6 74LS32
-21 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
8809 0 0
2
43055.8 3
0
9 2-In AND~
219 1120 339 0 3 22
0 22 21 16
0
0 0 112 0
6 74LS08
-21 -24 21 -16
4 U18A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 22 0
1 U
5993 0 0
2
43055.8 2
0
9 2-In XOR~
219 1043 311 0 3 22
0 11 23 22
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 U16B
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
8654 0 0
2
43055.8 1
0
9 2-In XOR~
219 960 320 0 3 22
0 12 19 23
0
0 0 112 0
6 74LS86
-21 -24 21 -16
4 U16C
-8 -25 20 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
7223 0 0
2
43055.8 0
0
14 Logic Display~
6 1238 673 0 1 2
10 24
0
0 0 53856 0
6 100MEG
3 -16 45 -8
1 S
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3641 0 0
2
43055.8 7
0
8 3-In OR~
219 1205 694 0 4 22
0 16 26 25 24
0
0 0 112 0
4 4075
-14 -24 14 -16
4 U14A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 18 0
1 U
3104 0 0
2
43055.8 9
0
8 4-In OR~
219 1038 796 0 5 22
0 34 33 32 31 25
0
0 0 112 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
3296 0 0
2
43055.8 24
0
8 4-In OR~
219 1040 591 0 5 22
0 30 29 28 27 26
0
0 0 112 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
8534 0 0
2
43055.8 25
0
9 2-In AND~
219 936 887 0 3 22
0 42 37 31
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
949 0 0
2
43055.8 26
0
9 2-In AND~
219 937 829 0 3 22
0 43 2 32
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
3371 0 0
2
43055.8 27
0
9 2-In AND~
219 938 779 0 3 22
0 44 35 33
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
7311 0 0
2
43055.8 28
0
9 2-In AND~
219 940 729 0 3 22
0 45 36 34
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 12 0
1 U
3409 0 0
2
43055.8 29
0
9 2-In AND~
219 939 676 0 3 22
0 46 38 27
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
3526 0 0
2
43055.8 30
0
9 2-In AND~
219 938 622 0 3 22
0 47 39 28
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 6 0
1 U
4129 0 0
2
43055.8 31
0
9 2-In AND~
219 937 570 0 3 22
0 48 40 29
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 6 0
1 U
6278 0 0
2
43055.8 32
0
9 2-In AND~
219 936 518 0 3 22
0 49 41 30
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
3482 0 0
2
43055.8 33
0
9 Inverter~
13 880 896 0 2 22
0 11 37
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U1F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 1 0
1 U
8323 0 0
2
43055.8 34
0
6 74266~
219 865 837 0 3 22
0 11 12 2
0
0 0 112 0
7 74LS266
-24 -24 25 -16
3 U7A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3984 0 0
2
43055.8 35
0
6 74136~
219 876 787 0 3 22
0 11 12 35
0
0 0 112 0
7 74LS136
-24 -24 25 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
7622 0 0
2
43055.8 36
0
9 2-In NOR~
219 875 737 0 3 22
0 58 12 36
0
0 0 112 0
6 74LS02
-21 -24 21 -16
3 U5A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 512 4 1 9 0
1 U
816 0 0
2
43055.8 37
0
8 2-In OR~
219 875 685 0 3 22
0 11 12 38
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 8 0
1 U
4656 0 0
2
43055.8 38
0
10 2-In NAND~
219 886 631 0 3 22
0 11 12 39
0
0 0 112 0
4 7400
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
6356 0 0
2
43055.8 39
0
9 2-In AND~
219 885 578 0 3 22
0 11 12 40
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
7479 0 0
2
43055.8 40
0
9 Inverter~
13 880 527 0 2 22
0 12 41
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U1E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 1 0
1 U
5690 0 0
2
43055.8 41
0
9 4-In AND~
219 746 879 0 5 22
0 50 54 52 57 42
0
0 0 624 0
3 NOT
-11 -28 10 -20
3 NOT
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
5617 0 0
2
43055.8 42
0
9 4-In AND~
219 746 823 0 5 22
0 53 51 55 57 43
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 XNOR
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
3903 0 0
2
43055.8 43
0
9 4-In AND~
219 745 772 0 5 22
0 56 52 54 50 44
0
0 0 624 0
6 74LS21
-21 -28 21 -20
3 XOR
-12 -28 9 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 2 0
1 U
4452 0 0
2
43055.8 44
0
5 7415~
219 743 667 0 4 22
0 52 51 50 46
0
0 0 624 0
6 74LS15
-21 -28 21 -20
2 OR
-9 -25 5 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 4 0
1 U
6282 0 0
2
43055.8 45
0
5 7415~
219 743 720 0 4 22
0 52 54 53 45
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 NOR
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 4 0
1 U
7187 0 0
2
43055.8 46
0
5 7415~
219 744 614 0 4 22
0 52 51 53 47
0
0 0 624 0
6 74LS15
-21 -28 21 -20
4 NAND
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 4 0
1 U
6866 0 0
2
43055.8 47
0
5 7415~
219 744 561 0 4 22
0 55 54 50 48
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 3 0
1 U
7670 0 0
2
43055.8 48
0
5 7415~
219 743 509 0 4 22
0 55 54 53 49
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 NOT
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 3 0
1 U
951 0 0
2
43055.8 49
0
5 7415~
219 742 394 0 4 22
0 55 51 50 7
0
0 0 624 0
6 74LS15
-21 -28 21 -20
3 SUB
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 3 0
1 U
9536 0 0
2
43055.8 50
0
9 4-In AND~
219 742 339 0 5 22
0 56 55 51 53 5
0
0 0 624 0
6 74LS21
-21 -28 21 -20
4 SOMA
-15 -28 13 -20
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 2 0
1 U
5495 0 0
2
43055.8 51
0
9 Inverter~
13 677 258 0 2 22
0 50 53
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
8152 0 0
2
43055.8 52
0
9 Inverter~
13 618 260 0 2 22
0 54 51
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
6223 0 0
2
43055.8 53
0
9 Inverter~
13 556 259 0 2 22
0 52 55
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
5441 0 0
2
43055.8 54
0
9 Inverter~
13 486 260 0 2 22
0 57 56
0
0 0 112 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
3189 0 0
2
43055.8 55
0
110
3 2 2 0 0 8320 0 36 28 0 0 3
904 837
904 838
913 838
1 3 3 0 0 0 0 8 9 0 0 2
1211 432
1211 432
3 1 4 0 0 8320 0 17 15 0 0 4
936 413
946 413
946 429
954 429
0 1 5 0 0 8192 0 0 17 27 0 3
790 339
790 404
891 404
3 1 6 0 0 8320 0 15 13 0 0 3
1003 438
1016 438
1016 468
1 4 7 0 0 4096 0 16 51 0 0 3
890 449
763 449
763 394
2 0 7 0 0 12288 0 10 0 0 8 4
1092 410
971 410
971 377
763 377
2 4 7 0 0 4224 0 19 51 0 0 3
987 357
763 357
763 394
1 3 8 0 0 8320 0 12 11 0 0 3
1094 459
1075 459
1075 374
3 2 9 0 0 4224 0 13 12 0 0 2
1061 477
1094 477
3 2 10 0 0 4224 0 14 13 0 0 2
1001 486
1016 486
0 1 5 0 0 0 0 0 19 27 0 2
955 339
987 339
1 0 11 0 0 4096 0 36 0 0 29 2
849 828
831 828
1 0 11 0 0 4096 0 37 0 0 29 2
860 778
831 778
1 0 11 0 0 4096 0 39 0 0 29 2
862 676
831 676
1 0 11 0 0 0 0 40 0 0 29 2
862 622
831 622
1 0 11 0 0 0 0 41 0 0 29 2
861 569
831 569
2 0 12 0 0 4096 0 40 0 0 28 2
862 640
853 640
2 0 12 0 0 0 0 41 0 0 28 2
861 587
853 587
1 0 12 0 0 4096 0 42 0 0 28 2
865 527
853 527
2 0 12 0 0 0 0 39 0 0 28 2
862 694
853 694
2 0 12 0 0 0 0 38 0 0 28 2
862 746
853 746
2 0 12 0 0 0 0 37 0 0 28 2
860 796
853 796
0 0 13 0 0 0 0 0 0 0 0 2
831 745
831 745
3 2 14 0 0 8320 0 12 9 0 0 4
1140 468
1156 468
1156 441
1166 441
3 1 15 0 0 8320 0 10 9 0 0 7
1138 401
1156 401
1156 423
1165 423
1165 424
1166 424
1166 423
5 1 5 0 0 4224 0 52 10 0 0 4
763 339
955 339
955 392
1092 392
1 2 12 0 0 4224 0 1 36 0 0 3
853 263
853 846
849 846
1 1 11 0 0 4224 0 2 35 0 0 3
831 263
831 896
865 896
1 0 11 0 0 0 0 2 0 0 0 2
831 263
831 504
3 1 16 0 0 8320 0 20 24 0 0 4
1141 339
1148 339
1148 685
1192 685
4 0 17 0 0 4224 0 0 0 0 0 2
764 339
843 339
1 2 11 0 0 0 0 2 17 0 0 3
831 263
831 422
891 422
2 2 18 0 0 4224 0 18 16 0 0 3
813 298
813 467
890 467
1 2 19 0 0 4224 0 3 14 0 0 3
880 264
880 495
955 495
1 1 12 0 0 0 0 1 14 0 0 3
853 263
853 477
955 477
1 2 19 0 0 0 0 3 11 0 0 3
880 264
880 383
1030 383
1 1 12 0 0 0 0 1 11 0 0 3
853 263
853 365
1030 365
3 2 20 0 0 8320 0 16 15 0 0 4
935 458
945 458
945 447
954 447
1 1 11 0 0 0 0 2 18 0 0 3
831 263
831 262
813 262
3 2 21 0 0 4224 0 19 20 0 0 2
1033 348
1096 348
3 1 22 0 0 8320 0 21 20 0 0 4
1076 311
1089 311
1089 330
1096 330
1 1 12 0 0 0 0 1 22 0 0 3
853 263
853 311
944 311
1 2 19 0 0 0 0 3 22 0 0 3
880 264
880 329
944 329
1 1 11 0 0 0 0 2 21 0 0 3
831 263
831 302
1027 302
3 2 23 0 0 4224 0 22 21 0 0 2
993 320
1027 320
1 4 24 0 0 8320 0 23 24 0 0 4
1238 691
1237 691
1237 694
1238 694
5 3 25 0 0 8320 0 25 24 0 0 4
1071 796
1135 796
1135 703
1192 703
5 2 26 0 0 8320 0 26 24 0 0 4
1073 591
1135 591
1135 694
1193 694
3 4 27 0 0 8320 0 31 26 0 0 4
960 676
980 676
980 605
1023 605
3 3 28 0 0 12416 0 32 26 0 0 4
959 622
971 622
971 596
1023 596
3 2 29 0 0 12416 0 33 26 0 0 4
958 570
971 570
971 587
1023 587
3 1 30 0 0 8320 0 34 26 0 0 4
957 518
980 518
980 578
1023 578
3 4 31 0 0 8320 0 27 25 0 0 4
957 887
980 887
980 810
1021 810
3 3 32 0 0 12416 0 28 25 0 0 4
958 829
972 829
972 801
1021 801
3 2 33 0 0 12416 0 29 25 0 0 4
959 779
972 779
972 792
1021 792
3 1 34 0 0 8320 0 30 25 0 0 4
961 729
980 729
980 783
1021 783
3 2 35 0 0 12416 0 37 29 0 0 4
909 787
906 787
906 788
914 788
3 2 36 0 0 4224 0 38 30 0 0 3
914 737
916 737
916 738
2 2 37 0 0 4224 0 35 27 0 0 2
901 896
912 896
3 2 38 0 0 4224 0 39 31 0 0 2
908 685
915 685
3 2 39 0 0 4224 0 40 32 0 0 2
913 631
914 631
3 2 40 0 0 8320 0 41 33 0 0 3
906 578
906 579
913 579
2 2 41 0 0 4224 0 42 34 0 0 2
901 527
912 527
5 1 42 0 0 8320 0 43 27 0 0 3
767 879
767 878
912 878
5 1 43 0 0 8320 0 44 28 0 0 3
767 823
767 820
913 820
5 1 44 0 0 8320 0 45 29 0 0 3
766 772
766 770
914 770
4 1 45 0 0 4224 0 47 30 0 0 2
764 720
916 720
4 1 46 0 0 4224 0 46 31 0 0 2
764 667
915 667
4 1 47 0 0 8320 0 48 32 0 0 3
765 614
765 613
914 613
4 1 48 0 0 4224 0 49 33 0 0 2
765 561
913 561
4 1 49 0 0 4224 0 50 34 0 0 2
764 509
912 509
3 0 50 0 0 4096 0 46 0 0 106 2
719 676
654 676
2 0 51 0 0 4096 0 46 0 0 100 2
719 667
621 667
1 0 52 0 0 4096 0 46 0 0 108 2
719 658
536 658
3 0 53 0 0 4096 0 48 0 0 99 2
720 623
680 623
2 0 51 0 0 4096 0 48 0 0 100 2
720 614
621 614
1 0 52 0 0 4096 0 48 0 0 108 2
720 605
536 605
3 0 50 0 0 4096 0 49 0 0 106 2
720 570
654 570
2 0 54 0 0 4096 0 49 0 0 107 2
720 561
590 561
1 0 55 0 0 4096 0 49 0 0 101 2
720 552
559 552
1 0 52 0 0 0 0 47 0 0 108 2
719 711
536 711
2 0 54 0 0 0 0 47 0 0 107 2
719 720
590 720
3 0 53 0 0 0 0 47 0 0 99 2
719 729
680 729
3 0 53 0 0 0 0 50 0 0 99 2
719 518
680 518
2 0 54 0 0 0 0 50 0 0 107 2
719 509
590 509
1 0 55 0 0 0 0 50 0 0 101 2
719 500
559 500
3 0 50 0 0 0 0 51 0 0 106 2
718 403
654 403
2 0 51 0 0 0 0 51 0 0 100 2
718 394
621 394
1 0 55 0 0 0 0 51 0 0 101 2
718 385
559 385
4 0 53 0 0 0 0 52 0 0 99 2
718 353
680 353
3 0 51 0 0 0 0 52 0 0 100 2
718 344
621 344
2 0 55 0 0 0 0 52 0 0 101 2
718 335
559 335
1 0 56 0 0 4096 0 52 0 0 95 2
718 326
489 326
2 1 56 0 0 4224 0 56 45 0 0 3
489 278
489 759
721 759
2 0 52 0 0 4096 0 45 0 0 108 2
721 768
536 768
3 0 54 0 0 4096 0 45 0 0 107 2
721 777
590 777
4 0 50 0 0 4096 0 45 0 0 106 2
721 786
654 786
2 1 53 0 0 4224 0 53 44 0 0 3
680 276
680 810
722 810
2 2 51 0 0 4224 0 54 44 0 0 3
621 278
621 819
722 819
2 3 55 0 0 4224 0 55 44 0 0 3
559 277
559 828
722 828
0 1 50 0 0 0 0 0 53 106 0 3
654 225
680 225
680 240
0 1 54 0 0 0 0 0 54 107 0 3
590 230
621 230
621 242
0 1 52 0 0 0 0 0 55 108 0 3
536 229
559 229
559 241
4 0 57 0 0 4096 0 44 0 0 110 2
722 837
464 837
1 1 50 0 0 4224 0 4 43 0 0 3
654 222
654 866
722 866
1 2 54 0 0 4224 0 7 43 0 0 3
590 224
590 875
722 875
1 3 52 0 0 4224 0 6 43 0 0 3
536 224
536 884
722 884
1 1 57 0 0 0 0 5 56 0 0 3
464 223
489 223
489 242
1 4 57 0 0 4224 0 5 43 0 0 3
464 223
464 893
722 893
0
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
